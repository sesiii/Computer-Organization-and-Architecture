module xor_gate(input [3:0]a,b,output [3:0]result);
assign result=(a^b);
endmodule